
module clk_div4(
input clk_4Hz,
input sys_rsn,
output reg clk_1Hz
);
reg [2:0] cnt4;

always @(posedge clk_4Hz or negedge sys_rsn) begin
	if(!sys_rsn)
		cnt4<=2'b0;
	else 
		cnt4<=cnt4+2'b1;
end


always @(posedge clk_4Hz ) begin
	if(cnt4<=2'd3)
		clk_1Hz<=1'b0;
	else 
		clk_1Hz<=1'b1;
end

endmodule
